----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    14:15:14 10/25/2023 
-- Design Name: 
-- Module Name:    ddf - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity ddf is
    Port ( input : in  STD_LOGIC;
           clk : in  STD_LOGIC;
           rst : in  STD_LOGIC;
           output : out  STD_LOGIC);
end ddf;

architecture Behavioral of ddf is

signal sig_betw : STD_LOGIC;

begin

	p: process(clk, rst) begin
        if (rst = '1') then
           sig_betw <= '0';
           output <= '0';
		elsif rising_edge(clk) then
			sig_betw <= input;
			output <= sig_betw;
		end if;
	end process;
 
end Behavioral;
